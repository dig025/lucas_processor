// Create Date:    2018.10.15
// Module Name:    ALU 
// Project Name:   CSE141L
//
// Revision 2018.01.27
// Additional Comments: 
//   combinational (unclocked) ALU 
import definitions::*;			           // includes package "definitions"
module ALU(
  input        [7:0] InputA,             // data inputs
                     InputB,
  input        [2:0] OP,		           // ALU opcode, part of microcode
  output logic [7:0] Out,		           // or:  output reg [7:0] OUT,
  output logic       Zero                // output = zero flag
    );								    
	 
  op_mne op_mnemonic;			           // type enum: used for convenient waveform viewing
  
  always_comb begin
    Out = 0;                             // No Op = default
    case(OP)
      kADD : Out = InputA + InputB;      // add 
      kLSH : Out = InputA << 1;  	     // shift left 
		kRSH : Out = {1'b0, InputA[7:1]};  // shift right
		kXOR : Out = InputA ^ InputB;      // exclusive OR
      kAND : Out = InputA & InputB;      // bitwise AND
    endcase
  end

  always_comb							  // assign Zero = !Out;
    case(Out)
      'b0     : Zero = 1'b1;
	  default : Zero = 1'b0;
    endcase

  always_comb
    op_mnemonic = op_mne'(OP);			 // displays operation name in waveform viewer

endmodule